`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:39:57 09/28/2016 
// Design Name: 
// Module Name:    cwalk_fsm 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module cwalk_fsm(
    input clk,
    input reset,
    input c7,
    input tc,
    output walk,
    output hand,
    output num_on,
    output en
    );
	 
	 // You may change the I/O signals above if you don't need certain outputs, etc.

endmodule
